// srlcsAdder_tb.v
// Vincent Li
// 3/26/2019
`timescale 1ns / 1ps

module srlcsAdder_tb;


endmodule
